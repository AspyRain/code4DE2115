
module demo2_waterled (
	clk_clk,
	reset_reset_n,
	led_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	led_export;
endmodule
